library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;

entity IM is
    Port ( Address : in  STD_LOGIC_VECTOR (31 downto 0);
           Reset : in  STD_LOGIC;
           Instruction : out  STD_LOGIC_VECTOR (31 downto 0));
end IM;

architecture Arqim of IM is

type rom_type is array (63 downto 0) of std_logic_vector (31 downto 0);
signal ROM : rom_type := (	"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", 
									"00000000000000000000000000000000", 
									"00000001000000000000000000000000",
									"01111111111111111111111111101000", 
									"10100110000100000010000000000110",
									"10100100000100000010000000001111", 
									"00000001000000000000000000000000",
									"10000011110000111110000000000000", 
									"10010000000100000000000000010000",
									"00000001000000000000000000000000",
									"00000110101111111111111111110100", 
									"10000000101001000100000000010011",
									"00000001000000000000000000000000",
									"00000001000000000000000000000000",
									"00000001000000000000000000000000",
									"10100010000100000000000000010100",
									"00000001000000000000000000000000",
									"00000001000000000000000000000000",
									"10101000000001000110000000000001",
									"10100000000100000000000000010100",
									"00000001000000000000000000000000",
									"00000001000000000000000000000000",
									"10101000000001000000000000010010",
									"00000001000000000000000000000000",
									"00110110100000000000000000010000",
									"10000000101001000100000000010011",	
									"10100010000100000010000000000000",
									"10100000000100000010000000000000");

begin

    process (Reset,Address,rom)
    begin
        if (Reset='1') then
				Instruction <= "00000000000000000000000000000000";
		  else
            Instruction <= ROM(conv_integer(Address(5 downto 0)));  
        end if;
    end process;
end Arqim;

