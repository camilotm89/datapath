library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity mux_wm_rf is
    Port ( a : in  STD_LOGIC_VECTOR (5 downto 0);
           b : in  STD_LOGIC_VECTOR (5 downto 0);
           sel : in  STD_LOGIC;
           out_mux : out  STD_LOGIC_VECTOR (5 downto 0));
end mux_wm_rf;

architecture Behavioral of mux_wm_rf is

begin
	process(a,b,sel)
	begin
		if (sel = '0')then
			out_mux <= a;
		else
			out_mux <= b;
		end if;
	end process;

end Behavioral;